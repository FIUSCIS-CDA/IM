
///////////////////////////////////////////////////////////////////////////////////
// Testbench for Component: IM
// Package: FIUSCIS-CDA
// Course: CDA3102 (Computer Architecture), Florida International University
// Developer: Trevor Cickovski
// License: MIT, (C) 2020 All Rights Reserved
///////////////////////////////////////////////////////////////////////////////////


module testbench();
`include "../Test/Test.v"

///////////////////////////////////////////////////////////////////////////////////
// Input: addr (32-bit)
reg[31:0] addr;
///////////////////////////////////////////////////////////////////////////////////

///////////////////////////////////////////////////////////////////////////////////
// Output: data (32-bit)
wire[31:0] data;
///////////////////////////////////////////////////////////////////////////////////

IM IMemory(.a(addr), 
           .d(data));


initial begin
/////////////////////////////////////////////////////////////////////////////
// Populate with program data
$readmemh("instmem.dat",IMemory.memory);
/////////////////////////////////////////////////////////////////////////////
// Test: addr=8
addr=8;  #100; 
$display("Testing with addr=8: "); 
verifyEqual32(data, 32'b10001100000011110000000001000000);
$display("All tests passed.");
end

endmodule